module Inverter( A,nA);
 input A;
 output nA;
  not inv1(nA,A);
endmodule

// Simulation parameters
// A CLK 10 10
